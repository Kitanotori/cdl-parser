test0
test1.@a
test2.@a.@b
test3(x>y)
test4(x>y).@a
test5(x>y).@a.@b
"test6"
"test7".@a
"test8".@a.@b
"test9.@a".@b
"test10,	137-145:1H
test11(icl	<	uw)
test12(icl>uw1(agt>uw2,obj>uw3),icl>uw4).@attr1.@attr2
test13..
test14..@attr
"test15..".@attr
"test16.@attr".@attr
"test17..().@"(icl>uw).@attr
test18(icl>uw(agt>uw2,obj>uw3),icl>uw4(agt>uw5))
test19(icl< uw)
test20(icl	<uw)