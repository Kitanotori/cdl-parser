<01:"test1".@attr>
<02:test2.@attr1.@attr2>
<03:"">
<04:2>
<05:>
<06:16(10)>
