test0
test1.@attr
"test2"
"test3".@attr
test4..
test5..@attr
"test6..".@attr
"test7.@attr".@attr
test8(icl>uw)
test9(icl>uw).@attr
"test10..().@"(icl>uw).@attr
test11(icl>uw(agt>uw2,obj>uw3),icl>uw4(agt>uw5))
test12(icl>uw1(agt>uw2,obj>uw3),icl>uw4).@attr1.@attr2
test13(agt>thing,obj>role>effect)
test14(icl< uw)
.@test15,	137-145:1H
>1.@topic
