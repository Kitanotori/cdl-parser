<01:"test1".@attr>
<02:test2.@attr1.@attr2>
<03:"">
<04:2>
<05:>
<06:16(x>y)>
<07:16(x>y).@c>
<08:16(x>y).@c.@d>
<09:a(b>c(d>e,f<g)).@h.@i>