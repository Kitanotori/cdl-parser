{#
	<01:a(x s<y(h>i),k<l).@a1>
	{#02
		<2A:b>
		<2B:c>
		[2A d 2B]
	}
	[01 e 02]
}