[1 agt 2]
