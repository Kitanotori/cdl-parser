<01:"test1".@attr>
<02:test2.@attr1.@attr2>
<03:"">
<04:2>
<05:>
<06:16(x>y)>
<07:16(x>y).@c>
<08:16(x>y).@c.@d>
<09:a(b>c(d>e,f<g)).@h.@i>
<10:a b.@c>
<11:3.0>
<12:3.0.@a>
<13:3.0(a>b).@c>
<14:etc.>
<15:etc..@a>
<16:etc.(a>b).@c>